-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : ALU
-- Author      : Judah Ben-Eliezer
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\SIMD\ALU\compile\SLIMAHS.vhd
-- Generated   : Sun Mar 28 22:23:34 2021
-- From        : C:\My_Designs\SIMD\ALU\..\blocks\SLIMAHS.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library ieee;
use ieee.std_logic_1164.all;
use ieee.NUMERIC_STD.all;

entity SLIMAHS is
  port(
       op : in STD_LOGIC_VECTOR(24 downto 0);
       i : in STD_LOGIC_VECTOR(127 downto 0);
       j : in STD_LOGIC_VECTOR(127 downto 0);
       k : in STD_LOGIC_VECTOR(127 downto 0);
       r : out STD_LOGIC_VECTOR(127 downto 0)
  );
end SLIMAHS;

architecture behavioral of SLIMAHS is

---- Component declarations -----

component MULT_ADD_L
  port(
       x : in STD_LOGIC_VECTOR(31 downto 0);
       y : in STD_LOGIC_VECTOR(31 downto 0);
       z : in STD_LOGIC_VECTOR(63 downto 0);
       result : out STD_LOGIC_VECTOR(63 downto 0)
  );
end component;

---- Signal declarations used on the diagram ----

signal res : STD_LOGIC_VECTOR(127 downto 0);

begin

---- Processes ----

process (op)
                       begin
                         if (op(24 downto 20) = "10101") then
                            r <= res;
                         end if;
                       end process;
                      

----  Component instantiations  ----

SLIMAHS_0 : MULT_ADD_L
  port map(
       x(31) => i(63),
       x(30) => i(62),
       x(29) => i(61),
       x(28) => i(60),
       x(27) => i(59),
       x(26) => i(58),
       x(25) => i(57),
       x(24) => i(56),
       x(23) => i(55),
       x(22) => i(54),
       x(21) => i(53),
       x(20) => i(52),
       x(19) => i(51),
       x(18) => i(50),
       x(17) => i(49),
       x(16) => i(48),
       x(15) => i(47),
       x(14) => i(46),
       x(13) => i(45),
       x(12) => i(44),
       x(11) => i(43),
       x(10) => i(42),
       x(9) => i(41),
       x(8) => i(40),
       x(7) => i(39),
       x(6) => i(38),
       x(5) => i(37),
       x(4) => i(36),
       x(3) => i(35),
       x(2) => i(34),
       x(1) => i(33),
       x(0) => i(32),
       y(31) => j(63),
       y(30) => j(62),
       y(29) => j(61),
       y(28) => j(60),
       y(27) => j(59),
       y(26) => j(58),
       y(25) => j(57),
       y(24) => j(56),
       y(23) => j(55),
       y(22) => j(54),
       y(21) => j(53),
       y(20) => j(52),
       y(19) => j(51),
       y(18) => j(50),
       y(17) => j(49),
       y(16) => j(48),
       y(15) => j(47),
       y(14) => j(46),
       y(13) => j(45),
       y(12) => j(44),
       y(11) => j(43),
       y(10) => j(42),
       y(9) => j(41),
       y(8) => j(40),
       y(7) => j(39),
       y(6) => j(38),
       y(5) => j(37),
       y(4) => j(36),
       y(3) => j(35),
       y(2) => j(34),
       y(1) => j(33),
       y(0) => j(32),
       z(63) => k(63),
       z(62) => k(62),
       z(61) => k(61),
       z(60) => k(60),
       z(59) => k(59),
       z(58) => k(58),
       z(57) => k(57),
       z(56) => k(56),
       z(55) => k(55),
       z(54) => k(54),
       z(53) => k(53),
       z(52) => k(52),
       z(51) => k(51),
       z(50) => k(50),
       z(49) => k(49),
       z(48) => k(48),
       z(47) => k(47),
       z(46) => k(46),
       z(45) => k(45),
       z(44) => k(44),
       z(43) => k(43),
       z(42) => k(42),
       z(41) => k(41),
       z(40) => k(40),
       z(39) => k(39),
       z(38) => k(38),
       z(37) => k(37),
       z(36) => k(36),
       z(35) => k(35),
       z(34) => k(34),
       z(33) => k(33),
       z(32) => k(32),
       z(31) => k(31),
       z(30) => k(30),
       z(29) => k(29),
       z(28) => k(28),
       z(27) => k(27),
       z(26) => k(26),
       z(25) => k(25),
       z(24) => k(24),
       z(23) => k(23),
       z(22) => k(22),
       z(21) => k(21),
       z(20) => k(20),
       z(19) => k(19),
       z(18) => k(18),
       z(17) => k(17),
       z(16) => k(16),
       z(15) => k(15),
       z(14) => k(14),
       z(13) => k(13),
       z(12) => k(12),
       z(11) => k(11),
       z(10) => k(10),
       z(9) => k(9),
       z(8) => k(8),
       z(7) => k(7),
       z(6) => k(6),
       z(5) => k(5),
       z(4) => k(4),
       z(3) => k(3),
       z(2) => k(2),
       z(1) => k(1),
       z(0) => k(0),
       result(63) => res(63),
       result(62) => res(62),
       result(61) => res(61),
       result(60) => res(60),
       result(59) => res(59),
       result(58) => res(58),
       result(57) => res(57),
       result(56) => res(56),
       result(55) => res(55),
       result(54) => res(54),
       result(53) => res(53),
       result(52) => res(52),
       result(51) => res(51),
       result(50) => res(50),
       result(49) => res(49),
       result(48) => res(48),
       result(47) => res(47),
       result(46) => res(46),
       result(45) => res(45),
       result(44) => res(44),
       result(43) => res(43),
       result(42) => res(42),
       result(41) => res(41),
       result(40) => res(40),
       result(39) => res(39),
       result(38) => res(38),
       result(37) => res(37),
       result(36) => res(36),
       result(35) => res(35),
       result(34) => res(34),
       result(33) => res(33),
       result(32) => res(32),
       result(31) => res(31),
       result(30) => res(30),
       result(29) => res(29),
       result(28) => res(28),
       result(27) => res(27),
       result(26) => res(26),
       result(25) => res(25),
       result(24) => res(24),
       result(23) => res(23),
       result(22) => res(22),
       result(21) => res(21),
       result(20) => res(20),
       result(19) => res(19),
       result(18) => res(18),
       result(17) => res(17),
       result(16) => res(16),
       result(15) => res(15),
       result(14) => res(14),
       result(13) => res(13),
       result(12) => res(12),
       result(11) => res(11),
       result(10) => res(10),
       result(9) => res(9),
       result(8) => res(8),
       result(7) => res(7),
       result(6) => res(6),
       result(5) => res(5),
       result(4) => res(4),
       result(3) => res(3),
       result(2) => res(2),
       result(1) => res(1),
       result(0) => res(0)
  );

SLIMAHS_1 : MULT_ADD_L
  port map(
       x(31) => i(127),
       x(30) => i(126),
       x(29) => i(125),
       x(28) => i(124),
       x(27) => i(123),
       x(26) => i(122),
       x(25) => i(121),
       x(24) => i(120),
       x(23) => i(119),
       x(22) => i(118),
       x(21) => i(117),
       x(20) => i(116),
       x(19) => i(115),
       x(18) => i(114),
       x(17) => i(113),
       x(16) => i(112),
       x(15) => i(111),
       x(14) => i(110),
       x(13) => i(109),
       x(12) => i(108),
       x(11) => i(107),
       x(10) => i(106),
       x(9) => i(105),
       x(8) => i(104),
       x(7) => i(103),
       x(6) => i(102),
       x(5) => i(101),
       x(4) => i(100),
       x(3) => i(99),
       x(2) => i(98),
       x(1) => i(97),
       x(0) => i(96),
       y(31) => j(127),
       y(30) => j(126),
       y(29) => j(125),
       y(28) => j(124),
       y(27) => j(123),
       y(26) => j(122),
       y(25) => j(121),
       y(24) => j(120),
       y(23) => j(119),
       y(22) => j(118),
       y(21) => j(117),
       y(20) => j(116),
       y(19) => j(115),
       y(18) => j(114),
       y(17) => j(113),
       y(16) => j(112),
       y(15) => j(111),
       y(14) => j(110),
       y(13) => j(109),
       y(12) => j(108),
       y(11) => j(107),
       y(10) => j(106),
       y(9) => j(105),
       y(8) => j(104),
       y(7) => j(103),
       y(6) => j(102),
       y(5) => j(101),
       y(4) => j(100),
       y(3) => j(99),
       y(2) => j(98),
       y(1) => j(97),
       y(0) => j(96),
       z(63) => k(127),
       z(62) => k(126),
       z(61) => k(125),
       z(60) => k(124),
       z(59) => k(123),
       z(58) => k(122),
       z(57) => k(121),
       z(56) => k(120),
       z(55) => k(119),
       z(54) => k(118),
       z(53) => k(117),
       z(52) => k(116),
       z(51) => k(115),
       z(50) => k(114),
       z(49) => k(113),
       z(48) => k(112),
       z(47) => k(111),
       z(46) => k(110),
       z(45) => k(109),
       z(44) => k(108),
       z(43) => k(107),
       z(42) => k(106),
       z(41) => k(105),
       z(40) => k(104),
       z(39) => k(103),
       z(38) => k(102),
       z(37) => k(101),
       z(36) => k(100),
       z(35) => k(99),
       z(34) => k(98),
       z(33) => k(97),
       z(32) => k(96),
       z(31) => k(95),
       z(30) => k(94),
       z(29) => k(93),
       z(28) => k(92),
       z(27) => k(91),
       z(26) => k(90),
       z(25) => k(89),
       z(24) => k(88),
       z(23) => k(87),
       z(22) => k(86),
       z(21) => k(85),
       z(20) => k(84),
       z(19) => k(83),
       z(18) => k(82),
       z(17) => k(81),
       z(16) => k(80),
       z(15) => k(79),
       z(14) => k(78),
       z(13) => k(77),
       z(12) => k(76),
       z(11) => k(75),
       z(10) => k(74),
       z(9) => k(73),
       z(8) => k(72),
       z(7) => k(71),
       z(6) => k(70),
       z(5) => k(69),
       z(4) => k(68),
       z(3) => k(67),
       z(2) => k(66),
       z(1) => k(65),
       z(0) => k(64),
       result(63) => res(127),
       result(62) => res(126),
       result(61) => res(125),
       result(60) => res(124),
       result(59) => res(123),
       result(58) => res(122),
       result(57) => res(121),
       result(56) => res(120),
       result(55) => res(119),
       result(54) => res(118),
       result(53) => res(117),
       result(52) => res(116),
       result(51) => res(115),
       result(50) => res(114),
       result(49) => res(113),
       result(48) => res(112),
       result(47) => res(111),
       result(46) => res(110),
       result(45) => res(109),
       result(44) => res(108),
       result(43) => res(107),
       result(42) => res(106),
       result(41) => res(105),
       result(40) => res(104),
       result(39) => res(103),
       result(38) => res(102),
       result(37) => res(101),
       result(36) => res(100),
       result(35) => res(99),
       result(34) => res(98),
       result(33) => res(97),
       result(32) => res(96),
       result(31) => res(95),
       result(30) => res(94),
       result(29) => res(93),
       result(28) => res(92),
       result(27) => res(91),
       result(26) => res(90),
       result(25) => res(89),
       result(24) => res(88),
       result(23) => res(87),
       result(22) => res(86),
       result(21) => res(85),
       result(20) => res(84),
       result(19) => res(83),
       result(18) => res(82),
       result(17) => res(81),
       result(16) => res(80),
       result(15) => res(79),
       result(14) => res(78),
       result(13) => res(77),
       result(12) => res(76),
       result(11) => res(75),
       result(10) => res(74),
       result(9) => res(73),
       result(8) => res(72),
       result(7) => res(71),
       result(6) => res(70),
       result(5) => res(69),
       result(4) => res(68),
       result(3) => res(67),
       result(2) => res(66),
       result(1) => res(65),
       result(0) => res(64)
  );


end behavioral;
