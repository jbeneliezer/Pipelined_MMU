-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : ALU
-- Author      : Judah Ben-Eliezer
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\SIMD\ALU\compile\SLIMALS.vhd
-- Generated   : Sun Mar 28 22:23:35 2021
-- From        : C:\My_Designs\SIMD\ALU\..\blocks\SLIMALS.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library ieee;
use ieee.std_logic_1164.all;
use ieee.NUMERIC_STD.all;

entity SLIMALS is
  port(
       op : in STD_LOGIC_VECTOR(24 downto 0);
       i : in STD_LOGIC_VECTOR(127 downto 0);
       j : in STD_LOGIC_VECTOR(127 downto 0);
       k : in STD_LOGIC_VECTOR(127 downto 0);
       r : out STD_LOGIC_VECTOR(127 downto 0)
  );
end SLIMALS;

architecture behavioral of SLIMALS is

---- Component declarations -----

component MULT_ADD_L
  port(
       x : in STD_LOGIC_VECTOR(31 downto 0);
       y : in STD_LOGIC_VECTOR(31 downto 0);
       z : in STD_LOGIC_VECTOR(63 downto 0);
       result : out STD_LOGIC_VECTOR(63 downto 0)
  );
end component;

---- Signal declarations used on the diagram ----

signal res : STD_LOGIC_VECTOR(127 downto 0);

begin

---- Processes ----

process (op)
                       begin
                         if (op(24 downto 20) = "10100") then
                            r <= res;
                         end if;
                       end process;
                      

----  Component instantiations  ----

SLIMALS_0 : MULT_ADD_L
  port map(
       x(31) => i(31),
       x(30) => i(30),
       x(29) => i(29),
       x(28) => i(28),
       x(27) => i(27),
       x(26) => i(26),
       x(25) => i(25),
       x(24) => i(24),
       x(23) => i(23),
       x(22) => i(22),
       x(21) => i(21),
       x(20) => i(20),
       x(19) => i(19),
       x(18) => i(18),
       x(17) => i(17),
       x(16) => i(16),
       x(15) => i(15),
       x(14) => i(14),
       x(13) => i(13),
       x(12) => i(12),
       x(11) => i(11),
       x(10) => i(10),
       x(9) => i(9),
       x(8) => i(8),
       x(7) => i(7),
       x(6) => i(6),
       x(5) => i(5),
       x(4) => i(4),
       x(3) => i(3),
       x(2) => i(2),
       x(1) => i(1),
       x(0) => i(0),
       y(31) => j(31),
       y(30) => j(30),
       y(29) => j(29),
       y(28) => j(28),
       y(27) => j(27),
       y(26) => j(26),
       y(25) => j(25),
       y(24) => j(24),
       y(23) => j(23),
       y(22) => j(22),
       y(21) => j(21),
       y(20) => j(20),
       y(19) => j(19),
       y(18) => j(18),
       y(17) => j(17),
       y(16) => j(16),
       y(15) => j(15),
       y(14) => j(14),
       y(13) => j(13),
       y(12) => j(12),
       y(11) => j(11),
       y(10) => j(10),
       y(9) => j(9),
       y(8) => j(8),
       y(7) => j(7),
       y(6) => j(6),
       y(5) => j(5),
       y(4) => j(4),
       y(3) => j(3),
       y(2) => j(2),
       y(1) => j(1),
       y(0) => j(0),
       z(63) => k(63),
       z(62) => k(62),
       z(61) => k(61),
       z(60) => k(60),
       z(59) => k(59),
       z(58) => k(58),
       z(57) => k(57),
       z(56) => k(56),
       z(55) => k(55),
       z(54) => k(54),
       z(53) => k(53),
       z(52) => k(52),
       z(51) => k(51),
       z(50) => k(50),
       z(49) => k(49),
       z(48) => k(48),
       z(47) => k(47),
       z(46) => k(46),
       z(45) => k(45),
       z(44) => k(44),
       z(43) => k(43),
       z(42) => k(42),
       z(41) => k(41),
       z(40) => k(40),
       z(39) => k(39),
       z(38) => k(38),
       z(37) => k(37),
       z(36) => k(36),
       z(35) => k(35),
       z(34) => k(34),
       z(33) => k(33),
       z(32) => k(32),
       z(31) => k(31),
       z(30) => k(30),
       z(29) => k(29),
       z(28) => k(28),
       z(27) => k(27),
       z(26) => k(26),
       z(25) => k(25),
       z(24) => k(24),
       z(23) => k(23),
       z(22) => k(22),
       z(21) => k(21),
       z(20) => k(20),
       z(19) => k(19),
       z(18) => k(18),
       z(17) => k(17),
       z(16) => k(16),
       z(15) => k(15),
       z(14) => k(14),
       z(13) => k(13),
       z(12) => k(12),
       z(11) => k(11),
       z(10) => k(10),
       z(9) => k(9),
       z(8) => k(8),
       z(7) => k(7),
       z(6) => k(6),
       z(5) => k(5),
       z(4) => k(4),
       z(3) => k(3),
       z(2) => k(2),
       z(1) => k(1),
       z(0) => k(0),
       result(63) => res(63),
       result(62) => res(62),
       result(61) => res(61),
       result(60) => res(60),
       result(59) => res(59),
       result(58) => res(58),
       result(57) => res(57),
       result(56) => res(56),
       result(55) => res(55),
       result(54) => res(54),
       result(53) => res(53),
       result(52) => res(52),
       result(51) => res(51),
       result(50) => res(50),
       result(49) => res(49),
       result(48) => res(48),
       result(47) => res(47),
       result(46) => res(46),
       result(45) => res(45),
       result(44) => res(44),
       result(43) => res(43),
       result(42) => res(42),
       result(41) => res(41),
       result(40) => res(40),
       result(39) => res(39),
       result(38) => res(38),
       result(37) => res(37),
       result(36) => res(36),
       result(35) => res(35),
       result(34) => res(34),
       result(33) => res(33),
       result(32) => res(32),
       result(31) => res(31),
       result(30) => res(30),
       result(29) => res(29),
       result(28) => res(28),
       result(27) => res(27),
       result(26) => res(26),
       result(25) => res(25),
       result(24) => res(24),
       result(23) => res(23),
       result(22) => res(22),
       result(21) => res(21),
       result(20) => res(20),
       result(19) => res(19),
       result(18) => res(18),
       result(17) => res(17),
       result(16) => res(16),
       result(15) => res(15),
       result(14) => res(14),
       result(13) => res(13),
       result(12) => res(12),
       result(11) => res(11),
       result(10) => res(10),
       result(9) => res(9),
       result(8) => res(8),
       result(7) => res(7),
       result(6) => res(6),
       result(5) => res(5),
       result(4) => res(4),
       result(3) => res(3),
       result(2) => res(2),
       result(1) => res(1),
       result(0) => res(0)
  );

SLIMALS_1 : MULT_ADD_L
  port map(
       x(31) => i(95),
       x(30) => i(94),
       x(29) => i(93),
       x(28) => i(92),
       x(27) => i(91),
       x(26) => i(90),
       x(25) => i(89),
       x(24) => i(88),
       x(23) => i(87),
       x(22) => i(86),
       x(21) => i(85),
       x(20) => i(84),
       x(19) => i(83),
       x(18) => i(82),
       x(17) => i(81),
       x(16) => i(80),
       x(15) => i(79),
       x(14) => i(78),
       x(13) => i(77),
       x(12) => i(76),
       x(11) => i(75),
       x(10) => i(74),
       x(9) => i(73),
       x(8) => i(72),
       x(7) => i(71),
       x(6) => i(70),
       x(5) => i(69),
       x(4) => i(68),
       x(3) => i(67),
       x(2) => i(66),
       x(1) => i(65),
       x(0) => i(64),
       y(31) => j(95),
       y(30) => j(94),
       y(29) => j(93),
       y(28) => j(92),
       y(27) => j(91),
       y(26) => j(90),
       y(25) => j(89),
       y(24) => j(88),
       y(23) => j(87),
       y(22) => j(86),
       y(21) => j(85),
       y(20) => j(84),
       y(19) => j(83),
       y(18) => j(82),
       y(17) => j(81),
       y(16) => j(80),
       y(15) => j(79),
       y(14) => j(78),
       y(13) => j(77),
       y(12) => j(76),
       y(11) => j(75),
       y(10) => j(74),
       y(9) => j(73),
       y(8) => j(72),
       y(7) => j(71),
       y(6) => j(70),
       y(5) => j(69),
       y(4) => j(68),
       y(3) => j(67),
       y(2) => j(66),
       y(1) => j(65),
       y(0) => j(64),
       z(63) => k(127),
       z(62) => k(126),
       z(61) => k(125),
       z(60) => k(124),
       z(59) => k(123),
       z(58) => k(122),
       z(57) => k(121),
       z(56) => k(120),
       z(55) => k(119),
       z(54) => k(118),
       z(53) => k(117),
       z(52) => k(116),
       z(51) => k(115),
       z(50) => k(114),
       z(49) => k(113),
       z(48) => k(112),
       z(47) => k(111),
       z(46) => k(110),
       z(45) => k(109),
       z(44) => k(108),
       z(43) => k(107),
       z(42) => k(106),
       z(41) => k(105),
       z(40) => k(104),
       z(39) => k(103),
       z(38) => k(102),
       z(37) => k(101),
       z(36) => k(100),
       z(35) => k(99),
       z(34) => k(98),
       z(33) => k(97),
       z(32) => k(96),
       z(31) => k(95),
       z(30) => k(94),
       z(29) => k(93),
       z(28) => k(92),
       z(27) => k(91),
       z(26) => k(90),
       z(25) => k(89),
       z(24) => k(88),
       z(23) => k(87),
       z(22) => k(86),
       z(21) => k(85),
       z(20) => k(84),
       z(19) => k(83),
       z(18) => k(82),
       z(17) => k(81),
       z(16) => k(80),
       z(15) => k(79),
       z(14) => k(78),
       z(13) => k(77),
       z(12) => k(76),
       z(11) => k(75),
       z(10) => k(74),
       z(9) => k(73),
       z(8) => k(72),
       z(7) => k(71),
       z(6) => k(70),
       z(5) => k(69),
       z(4) => k(68),
       z(3) => k(67),
       z(2) => k(66),
       z(1) => k(65),
       z(0) => k(64),
       result(63) => res(127),
       result(62) => res(126),
       result(61) => res(125),
       result(60) => res(124),
       result(59) => res(123),
       result(58) => res(122),
       result(57) => res(121),
       result(56) => res(120),
       result(55) => res(119),
       result(54) => res(118),
       result(53) => res(117),
       result(52) => res(116),
       result(51) => res(115),
       result(50) => res(114),
       result(49) => res(113),
       result(48) => res(112),
       result(47) => res(111),
       result(46) => res(110),
       result(45) => res(109),
       result(44) => res(108),
       result(43) => res(107),
       result(42) => res(106),
       result(41) => res(105),
       result(40) => res(104),
       result(39) => res(103),
       result(38) => res(102),
       result(37) => res(101),
       result(36) => res(100),
       result(35) => res(99),
       result(34) => res(98),
       result(33) => res(97),
       result(32) => res(96),
       result(31) => res(95),
       result(30) => res(94),
       result(29) => res(93),
       result(28) => res(92),
       result(27) => res(91),
       result(26) => res(90),
       result(25) => res(89),
       result(24) => res(88),
       result(23) => res(87),
       result(22) => res(86),
       result(21) => res(85),
       result(20) => res(84),
       result(19) => res(83),
       result(18) => res(82),
       result(17) => res(81),
       result(16) => res(80),
       result(15) => res(79),
       result(14) => res(78),
       result(13) => res(77),
       result(12) => res(76),
       result(11) => res(75),
       result(10) => res(74),
       result(9) => res(73),
       result(8) => res(72),
       result(7) => res(71),
       result(6) => res(70),
       result(5) => res(69),
       result(4) => res(68),
       result(3) => res(67),
       result(2) => res(66),
       result(1) => res(65),
       result(0) => res(64)
  );


end behavioral;
